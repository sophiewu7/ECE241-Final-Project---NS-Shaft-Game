		/*****************************************************************************
		 *                                                                           *
		 * Module:       Altera_UP_Audio_Bit_Counter                                 *
		 * Description:                                                              *
		 *      This module counts which bits for serial audio transfers. The module *
		 *   assume that the data format is I2S, as it is described in the audio     *
		 *   chip's datasheet.                                                       *
		 *                                                                           *
		 *****************************************************************************/

		module Altera_UP_Audio_Bit_Counter (
			// Inputs
			clk,
			reset,
			
			bit_clk_rising_edge,
			bit_clk_falling_edge,
			left_right_clk_rising_edge,
			left_right_clk_falling_edge,
			
			// Bidirectionals

			// Outputs
			counting
		);

		/*****************************************************************************
		 *                           Parameter Declarations                          *
		 *****************************************************************************/

		parameter BIT_COUNTER_INIT	= 5'd31;

		/*****************************************************************************
		 *                             Port Declarations                             *
		 *****************************************************************************/

		// Inputs
		input				clk;
		input				reset;
			
		input				bit_clk_rising_edge;
		input				bit_clk_falling_edge;
		input				left_right_clk_rising_edge;
		input				left_right_clk_falling_edge;

		// Bidirectionals

		// Outputs
		output	reg			counting;

		/*****************************************************************************
		 *                           Constant Declarations                           *
		 *****************************************************************************/


		/*****************************************************************************
		 *                 Internal wires and registers Declarations                 *
		 *****************************************************************************/

		// Internal Wires
		wire				reset_bit_counter;

		// Internal Registers
		reg			[4:0]	bit_counter;

		// State Machine Registers


		/*****************************************************************************
		 *                         Finite State Machine(s)                           *
		 *****************************************************************************/


		/*****************************************************************************
		 *                             Sequential logic                              *
		 *****************************************************************************/

		always @(posedge clk)
		begin
			if (reset == 1'b1)
				bit_counter <= 5'h00;
			else if (reset_bit_counter == 1'b1)
				bit_counter <= BIT_COUNTER_INIT;
			else if ((bit_clk_falling_edge == 1'b1) && (bit_counter != 5'h00))
				bit_counter <= bit_counter - 5'h01;
		end

		always @(posedge clk)
		begin
			if (reset == 1'b1)
				counting <= 1'b0;
			else if (reset_bit_counter == 1'b1)
				counting <= 1'b1;
			else if ((bit_clk_falling_edge == 1'b1) && (bit_counter == 5'h00))
				counting <= 1'b0;
		end

		/*****************************************************************************
		 *                            Combinational logic                            *
		 *****************************************************************************/

		assign reset_bit_counter = left_right_clk_rising_edge | 
									left_right_clk_falling_edge;

		/*****************************************************************************
		 *                              Internal Modules                             *
		 *****************************************************************************/

		endmodule

